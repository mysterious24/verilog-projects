module inv (a,out);
input a;
output out;

assign out=~a;
endmodule
